module SinglePulser (
    input syncpress_i,
    input clk, rst,
    output reg SP_o
);
    localparam S0 = 0, S1 = 1;
    reg state, next_state;

    always @(posedge clk) begin
        state <= (rst)? S0 : next_state;
    end

    always @* begin
        case (state)
            S0: begin
                next_state = (syncpress_i)? S1 : S0;
                SP_o = (syncpress_i)? 1 : 0;
            end
            S1: begin
                next_state = (syncpress_i)? S1 : S0;
                SP_o = 0;
            end
        endcase
    end
endmodule

module t_ShiftAddMultiplier (

);
endmodule
